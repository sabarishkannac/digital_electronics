`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/25/2025 11:31:03 AM
// Design Name: 
// Module Name: decoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module decoder( input [2:0] x ,output reg [7:0]  y);

always @(x)
begin
case(x)
3'b000:y=8'b00000000;
3'b001:y=8'b00000001;
3'b010:y=8'b00000010;
3'b011:y=8'b00000100;
3'b100:y=8'b00001000;
3'b101:y=8'b00010000;
3'b110:y=8'b00100000;
3'b111:y=8'b01000000;
endcase
end

endmodule
